module V1(clk,clk2,itemS,val,out,change,state);
input clk,clk2;
input [4:0] val,itemS;
output reg [4:0] state;
output reg [4:0]change;
output reg out;
parameter C0=0,C1=5,C2=10,C3=15,C4=20,C5=25,C6=30,C7=35,C8=40;
parameter none=0,Grape=1,Orange=2,Mango=3,Pineapple=4;
parameter S0=0,S1=1,S2=2,S3=3,S4=4,S5=5,S6=6,S7=7,S8=8;
always@(posedge clk)
begin 
    case(itemS)
    Grape:
    begin
        case(state)
        S0:
        begin
            if(val==5)
            state<=S1;
            else if(val==10)
            state<=S2;
            else if(val==20)
            state<=S4;
        end
        S1:
        begin 
            if(val==5)
            state<=S2;
            if(val==10)
            state<=S3;
            if(val==20)
            state<=S5;
        end
        S2:
        begin
            if(val==5)
            state<=S3;
            else if(val==10)
            state<=S4;
            else if(val==20)
            state<=S6;
        end
        S3:
        begin
            if(val==5)
            state<=S4;
            else if(val==10)
            state<=S5;
            else if(val==20)
            state<=S7;
        end
        S4:
        begin
            if(val==5)
            state<=S5;
            else if(val==10)
            state<=S6;
            else if(val==20)
            state<=S8;
        end
        S5:
        begin
            if(val==5)
            state<=S6;
            else if(val==10)
            state<=S7;
        end
        S6:
        if(val==5)
            state<=S7;
        else if(val==10)
            state<=S8;
        S7:
        if(val==5)
            state<=S8;
        S8:
        state<=S8;
        default:
        state<=S0;
    endcase
    end
    Orange:
    begin
        case(state)
        S0:
        begin
            if(val==5)
            state<=S1;
            else if(val==10)
            state<=S2;
            else if(val==20)
            state<=S4;
        end
        S1:
        begin 
            if(val==5)
            state<=S2;
            if(val==10)
            state<=S3;
            if(val==20)
            state<=S5;
        end
        S2:
        begin 
            if(val==5)
            state<=S3;
            if(val==10)
            state<=S4;
            if(val==20)
            state<=S6;
        end
        S3:
        begin
            if(val==5)
            state<=S4;
            else if(val==10)
            state<=S5;
            else if(val==20)
            state<=S7;
        end
        S4:
        begin
            if(val==5)
            state<=S5;
            else if(val==10)
            state<=S6;
            else if(val==20)
            state<=S8;
        end
        S5:
        begin
            if(val==5)
            state<=S6;
            else if(val==10)
            state<=S7;
        end
        S6:
        begin
            if(val==5)
            state<=S7;
            else if(val==10)
            state<=S8;
        end
        S7:
        begin
            if(val==5)
            state<=S8;
        end
        S8:
        state<=S8;
        default:
        state<=S0;
        endcase 
    end
    Mango:
    begin 
        case(state)
        S0:
        begin
            if(val==5)
            state<=S1;
            else if(val==10)
            state<=S2;
            else if(val==20)
            state<=S4;
        end
        S1:
        begin 
            if(val==5)
            state<=S2;
            if(val==10)
            state<=S3;
            if(val==20)
            state<=S5;
        end
        S2:
        begin 
            if(val==5)
            state<=S3;
            if(val==10)
            state<=S4;
            if(val==20)
            state<=S6;
        end
        S3:
        begin 
            if(val==5)
            state<=S4;
            if(val==10)
            state<=S5;
            if(val==20)
            state<=S7;
        end
        S4:
        begin
            if(val==5)
            state<=S5;
            else if(val==10)
            state<=S6;
            else if(val==20)
            state<=S8;
        end
        S5:
        begin
            if(val==5)
            state<=S6;
            else if(val==10)
            state<=S7;
        end
        S6:
        begin
            if(val==5)
            state<=S7;
            else if(val==10)
            state<=S8;
        end
        S7:
        begin
            if(val==5)
            state<=S8;
        end
        S8:
        state<=S8;
        default:
        state<=S0;
        endcase
    end
    Pineapple:
    begin
        case(state)
        S0:
        begin
            if(val==5)
            state<=S1;
            else if(val==10)
            state<=S2;
            else if(val==20)
            state<=S4;
        end
        S1:
        begin 
            if(val==5)
            state<=S2;
            if(val==10)
            state<=S3;
            if(val==20)
            state<=S5;
        end
        S2:
        begin 
            if(val==5)
            state<=S3;
            if(val==10)
            state<=S4;
            if(val==20)
            state<=S6;
        end
        S3:
        begin 
            if(val==5)
            state<=S4;
            if(val==10)
            state<=S5;
            if(val==20)
            state<=S7;
        end
        S4:
        begin 
            if(val==5)
            state<=S3;
            if(val==10)
            state<=S4;
            if(val==20)
            state<=S6;
        end
        S5:
        begin
            if(val==5)
            state<=S6;
            else if(val==10)
            state<=S7;
        end
        S6:
        begin
            if(val==5)
            state<=S7;
            else if(val==10)
            state<=S8;
        end
        S7:
        begin
            if(val==5)
            state<=S8;
        end
        S8:
        state<=S8;
        default:
        state<=S0;
        endcase
    end
    endcase
end
always@(posedge clk2)
begin 
    case(itemS)
    Grape:
        case(val)
        C1:
        begin 
            case(state)
                S0:begin
                out=0;change=0;end
                S1:begin
                out=1;change=0;end
                S2:begin
                out=1;change=5;end
                S3:begin
                out=1;change=10;end
                S4:begin
                out=1;change=15;end
                S5:begin
                out=1;change=20;end
                S6:begin
                out=1;change=25;end
                S7:begin
                out=5;change=30;end
            endcase
        end
        C2:
        begin 
            case(state)
                S0:begin
                out=1;change=0;end
                S1:begin
                out=1;change=5;end
                S2:begin
                out=1;change=10;end
                S3:begin
                out=1;change=15;end
                S4:begin
                out=1;change=20;end
                S5:begin
                out=1;change=25;end
                S6:begin
                out=1;change=30;end
                S7:begin
                out=5;change=35;end
            endcase
        end
        C4:
        begin 
            case(state)
                S0:begin
                out=1;change=10;end
                S1:begin
                out=1;change=15;end
                S2:begin
                out=1;change=20;end
                S3:begin
                out=1;change=25;end
                S4:begin
                out=1;change=30;end
                S5:begin
                out=1;change=40;end
                S6:begin
                out=1;change=45;end
                S7:begin
                out=5;change=50;end
            endcase
        end
        endcase
    Orange:
        case(val)
        C1:
        begin 
            case(state)
                S0:begin
                out=0;change=0;end
                S1:begin
                out=0;change=0;end
                S2:begin
                out=1;change=0;end
                S3:begin
                out=1;change=5;end
                S4:begin
                out=1;change=10;end
                S5:begin
                out=1;change=15;end
                S6:begin
                out=1;change=20;end
                S7:begin
                out=5;change=25;end
            endcase
        end
        C2:
        begin 
            case(state)
                S0:begin
                out=0;change=0;end
                S1:begin
                out=1;change=0;end
                S2:begin
                out=1;change=5;end
                S3:begin
                out=1;change=10;end
                S4:begin
                out=1;change=15;end
                S5:begin
                out=1;change=20;end
                S6:begin
                out=1;change=25;end
                S7:begin
                out=5;change=30;end
            endcase
        end
        C4:
        begin 
            case(state)
                S0:begin
                out=1;change=5;end
                S1:begin
                out=1;change=10;end
                S2:begin
                out=1;change=15;end
                S3:begin
                out=1;change=20;end
                S4:begin
                out=1;change=25;end
                S5:begin
                out=1;change=30;end
                S6:begin
                out=1;change=35;end
                S7:begin
                out=5;change=40;end
            endcase
        end
        endcase
    Mango:
        case(val)
        C1:
        begin 
            case(state)
                S0:begin
                out=0;change=0;end
                S1:begin
                out=0;change=0;end
                S2:begin
                out=0;change=0;end
                S3:begin
                out=1;change=0;end
                S4:begin
                out=1;change=5;end
                S5:begin
                out=1;change=10;end
                S6:begin
                out=1;change=15;end
                S7:begin
                out=5;change=20;end
            endcase
        end
        C2:
        begin 
            case(state)
                S0:begin
                out=0;change=0;end
                S1:begin
                out=0;change=0;end
                S2:begin
                out=1;change=0;end
                S3:begin
                out=1;change=5;end
                S4:begin
                out=1;change=10;end
                S5:begin
                out=1;change=15;end
                S6:begin
                out=1;change=20;end
                S7:begin
                out=5;change=25;end
            endcase
        end
        C4:
        begin 
            case(state)
                S0:begin
                out=1;change=0;end
                S1:begin
                out=1;change=5;end
                S2:begin
                out=1;change=10;end
                S3:begin
                out=1;change=15;end
                S4:begin
                out=1;change=20;end
                S5:begin
                out=1;change=25;end
                S6:begin
                out=1;change=30;end
                S7:begin
                out=1;change=35;end
            endcase
        end
        endcase
    Pineapple:
        case(val)
        C1:
        begin 
            case(state)
                S0:begin
                out=0;change=0;end
                S1:begin
                out=0;change=0;end
                S2:begin
                out=0;change=0;end
                S3:begin
                out=0;change=0;end
                S4:begin
                out=1;change=0;end
                S5:begin
                out=1;change=5;end
                S6:begin
                out=1;change=10;end
                S7:begin
                out=5;change=15;end
            endcase
        end
        C2:
        begin 
            case(state)
                S0:begin
                out=0;change=0;end
                S1:begin
                out=0;change=0;end
                S2:begin
                out=0;change=0;end
                S3:begin
                out=1;change=0;end
                S4:begin
                out=1;change=5;end
                S5:begin
                out=1;change=10;end
                S6:begin
                out=1;change=15;end
                S7:begin
                out=1;change=20;end
            endcase
        end
        C4:
        begin 
            case(state)
                S0:begin
                out=0;change=0;end
                S1:begin
                out=1;change=0;end
                S2:begin
                out=1;change=5;end
                S3:begin
                out=1;change=10;end
                S4:begin
                out=1;change=15;end
                S5:begin
                out=1;change=20;end
                S6:begin
                out=1;change=25;end
                S7:begin
                out=5;change=30;end
            endcase
        end
        endcase
    endcase
end
endmodule